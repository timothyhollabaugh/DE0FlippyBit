
module Column_State_Machine_Test()